`ifndef UTILS_PKG_SV
`define UTILS_PKG_SV

package utils_pkg;
	
endpackage : utils_pkg

`endif