package sum_pkg;
    import "DPI-C" function int add(int a, int b);
    import "DPI-C" function int getSum();
endpackage